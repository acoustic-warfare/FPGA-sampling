library IEEE;
use IEEE.STD_LOGIC_1164.all;

library vunit_lib;
context vunit_lib.vunit_context;

use work.MATRIX_TYPE.all;

entity tb_sample_clk is
   generic (
      runner_cfg : string
   );

end tb_sample_clk;

architecture behave of tb_sample_clk is
   constant C_CLK_CYKLE : time := 10 ns; -- set the duration of one clock cycle

   signal clk        : std_logic := '0';
   signal reset      : std_logic := '0';
   signal ws         : std_logic := '0';
   signal bit_stream : std_logic := '1';

   signal mic_sample_data_out  : std_logic_vector(23 downto 0);
   signal mic_sample_valid_out : std_logic;

   signal sim_counter : integer := 0;
   signal counter_tb  : integer := 0;

begin
   clk <= not(clk) after C_CLK_CYKLE/2;

   sample_clk1 : entity work.sample_clk
      generic map(
         index => 4
      )
      port map(
         sys_clk              => clk,
         reset                => reset,
         bit_stream           => bit_stream,
         ws                   => ws,
         mic_sample_data_out  => mic_sample_data_out,
         mic_sample_valid_out => mic_sample_valid_out
      );

   ws_process : process (clk)
   begin
      if falling_edge(clk) then
         if (counter_tb = 10 or counter_tb = 522*5 or counter_tb = 1034*5) then
            ws <= '1';
         else
            ws <= '0';
         end if;
         counter_tb <= counter_tb + 1;
      end if;
   end process;

   main : process
   begin
      test_runner_setup(runner, runner_cfg);
      while test_suite loop
         if run("wave") then
            -- test 1 is so far only ment for gktwave

            wait for 100000 ns; -- duration of test 1

         elsif run("auto") then

            wait for 11 ns;

         end if;
      end loop;

      test_runner_cleanup(runner);
   end process;

   test_runner_watchdog(runner, 100 ms);
end architecture;