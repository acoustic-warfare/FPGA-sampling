library ieee;
use ieee.std_logic_1164.all;

library vunit_lib;
context vunit_lib.vunit_context;

use work.matrix_type.all;

entity tb_clk_gen is
   generic (
      runner_cfg : string
   );
end tb_clk_gen;

architecture tb of tb_clk_gen is
   constant sck_cykle : time := 10 ns; -- set the duration of one clock cycle

   signal sck_clk : std_logic := '0';
   signal reset : std_logic;
   signal ws_pulse : std_logic;
   signal sck_counter : integer := 0; -- counter for the number of fsck_clk cycles
   signal ws_counter : integer := 0; -- counter for the number of fs_clk cykles

   signal auto : std_logic := '0';
   signal sck_counter_start : integer;

   procedure clk_wait (nr_of_cykles : in integer) is
   begin
      for i in 0 to nr_of_cykles loop
         wait for sck_cykle;
      end loop;
   end procedure;

begin
   -- direct instantiation of: clk_gen
   clk_gen_1 : entity work.clk_gen port map(
      sck_clk => sck_clk,
      ws_pulse => ws_pulse,
      reset => reset
      );

   -- counter for fs_clk cykles
   fsck_counter_p : process (sck_clk)
   begin
      if (rising_edge(sck_clk) and reset = '0') then
         sck_counter <= sck_counter + 1;
      end if;
   end process;

   -- counter for fs_clk cykles
   ws_counter_p : process (ws_pulse)
   begin
      if (rising_edge(ws_pulse) and reset = '0') then
         ws_counter <= ws_counter + 1;
      end if;
   end process;

   -- generate clock pulses with a clock period of clk_cykle
   clock_p : process
   begin
      sck_clk <= not(sck_clk);
      wait for sck_cykle/2;
   end process;

   assert_p : process (ws_pulse)
   begin
      if (auto = '1') then
         if (rising_edge(ws_pulse)) then
            if (ws_counter = 0) then
               sck_counter_start <= sck_counter;
            elsif (ws_counter = 1) then
               assert (sck_counter - sck_counter_start - 1 ) = 513 report "hej!" severity error; -- funkar inte rikgit �n
            end if;
         end if;
      end if;
   end process;

   main_p : process
   begin
      test_runner_setup(runner, runner_cfg);
      while test_suite loop
         if run("gkw") then -- only for use in gktwave

            reset <= '1';
            clk_wait(5);
            reset <= '0';

            wait for 30000 ns; -- duration of test 1

         elsif run("auto") then

            auto <= '1';
            reset <= '1';
            clk_wait(5);
            reset <= '0';

            wait for 100 ns; -- duration of test 1

         end if;
      end loop;

      test_runner_cleanup(runner);
   end process;

   test_runner_watchdog(runner, 100 ms);
end architecture;