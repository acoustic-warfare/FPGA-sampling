library ieee;
use ieee.std_logic_1164.all;
use work.matrix_type.all;
use ieee.numeric_std.all;
entity collector is
   ------------------------------------------------------------------------------------------------------------------------------------------------
   --                                                  # port information #
   -- MICID_SW: Signal to indicate if padding should be an ID for each mic or two's complement. 
   --
   -- MIC_SAMPLE_DATA_IN: Incomming array of data. One microphone sends 32 bits.
   --
   -- MIC_SAMPLE_VALID_IN: High for one clk cykle when the MIC_SAMPLE_DATA_IN has bean updated
   --
   -- CHAIN_MATRIX_DATA_OUT: A matrix filled the data from all the mics of the chain (16x32)
   --
   -- CHAIN_MATRIX_VALID_OUT: Indicates to the next component that the data has ben updated in CHAIN_MATRIX_DATA_OUT
   ------------------------------------------------------------------------------------------------------------------------------------------------
   generic (
      -- TODO: implement generics
      G_BITS_MIC : integer := 24; -- Defines the resulotion of a mic sample
      G_NR_MICS  : integer := 16; -- Number of chains in the Matrix
      chainID    : integer := 0   -- Identifier for a specific chain
   );
   port (
      sys_clk                : in std_logic;
      reset                  : in std_logic;
      micID_sw               : in std_logic;
      mic_sample_data_in     : in std_logic_vector(23 downto 0);
      mic_sample_valid_in    : in std_logic;
      chain_matrix_data_out  : out matrix_16_32_type; -- Our output Matrix with 1 sample from all microphones in the Matrix
      chain_matrix_valid_out : out std_logic := '0'   -- A signal to tell the receiver to start reading the data_out_matrix
   );
end collector;

architecture rtl of collector is
   signal counter_mic           : integer := 0; --Counter for rows in data_matrix_16_32_out
   signal mic_sample_valid_in_d : std_logic;
begin
   collect_p : process (sys_clk)                        -- Process which collects the input data and put it in the matrix
      variable tmp_holder : std_logic_vector(31 downto 0); -- temporary holder for incomming data, used for padding
   begin
      if rising_edge(sys_clk) then
         chain_matrix_valid_out <= '0';                                    -- Set data_valid_out to LOW as defult value
         if mic_sample_valid_in = '1' and mic_sample_valid_in_d = '0' then -- Data from a new mic is valid and the shift register puts it at the first place
            tmp_holder(23 downto 0) := mic_sample_data_in;
            if micID_sw = '0' then

               -- This part is not optimal but mabye necisary if we cant find a perfect delay :(
               if tmp_holder(23) = '1' and tmp_holder(22 downto 16) = "0000000" then
                  tmp_holder(23) := '0';
               elsif tmp_holder(23) = '0' and tmp_holder(22 downto 16) = "1111111" then
                  tmp_holder(23) := '1';
               elsif tmp_holder(22) = '1' and tmp_holder(21 downto 16) = "000000" then
                  tmp_holder(22) := '0';
               elsif tmp_holder(22) = '0' and tmp_holder(21 downto 16) = "111111" then
                  tmp_holder(22) := '1';
               end if;
               -- end of not optimal code

               if (tmp_holder(23) = '0') then
                  tmp_holder(31 downto 24) := "00000000"; -- Add padding according to TWO'S COMPLIMENT. if the 23:rd bit = 0 then padding = "00000000"
               else
                  tmp_holder(31 downto 24) := "11111111"; -- Add padding according to TWO'S COMPLIMENT. if the 23:rd bit = 1 then padding = "11111111"
               end if;
            else
               tmp_holder(31 downto 24) := std_logic_vector(to_unsigned(chainID * 16 + counter_mic, 8)); --Add padding according to the the current mic. if 2:nd mic then padding = "00000010"
            end if;

            chain_matrix_data_out(counter_mic) <= tmp_holder;
            counter_mic                        <= counter_mic + 1;
         end if;

         if counter_mic = 16 then -- When all Vectors is full in the matrix set the data_valid_out to HIGH
            chain_matrix_valid_out <= '1';
            counter_mic            <= 0; -- Resets the microphone counter, to prepare collect the chain again
         end if;

         mic_sample_valid_in_d <= mic_sample_valid_in;

         if reset = '1' then -- When reset is HIGH data_valid_out and counter_mic are reset back to LOW and zero
            chain_matrix_valid_out <= '0';
            counter_mic            <= 0;
         end if;
      end if;
   end process;
end rtl;